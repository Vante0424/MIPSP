
`include "define.v"
module InstMem(
    input wire ce,
    input wire [31:0] addr,
    output reg [31:0] data
);
    reg [31:0] instmem [1023 : 0];    
    always@(*)      
        if(ce == `RomDisable)
          data = `Zero;
        else
          data = instmem[addr[11 : 2]];   
    initial
      begin
	
		//ori
        instmem [0] = 32'h34011100;  //001101 00000 00001 0001000100000000  //ori r0 r1 1100
        instmem [1] = 32'h34020020;  //001101 00000 00010 0000000000100000  //ori r0 r2 0020
        instmem [2] = 32'h3403ff00;  //001101 00000 00011 1111111100000000  //ori r0 r3 ff00
        instmem [3] = 32'h3404ffff;  //001101 00000 00100 1111111111111111  //ori r0 r4 ffff
        
		//bgtz 6
		instmem [4] = 32'h1C200001;  //000111 00001 00000 0000000000000001  //bgtz r1
			
		//ori
		instmem [5] = 32'h34051100;  //001101 00000 00101 0001000100000000  //ori r0 r5 1100
		instmem [6] = 32'h34060028;  //001101 00000 00110 0000000000101000  //ori r0 r6 0028
		//slt (2 1 7)
		instmem [7] = 32'h0041382A;  //000000 00010 00001 00111 00000 101010  //slt r2 r1 r7
		//jalr 10(r6 zhuyi*4) cun 9 
		instmem [8] = 32'h00C0F809;  //000000 00110 00000 11111 00000 001001  //jalr 
		//ori 8 9 jicunqi 
		instmem [9] = 32'h34081100;   //001101 00000 01000 0001000100000000  //ori r0 r8 1100
		instmem [10] = 32'h34090020;  //001101 00000 01001 0000000000100000  //ori r0 r9 0020
		//multu r1 * r9 (un)
		instmem [11] = 32'h00290019;  //000000 00001 01001 00000 00000 011001  //multu r1 r9
		//hi -> r10
		instmem [12] = 32'h00005010;  //000000 00000 00000 01010 00000 010000  //mfhi r10
		//lo -> r11
		instmem [13] = 32'h00005812;  //000000 00000 00000 01011 00000 010010  //mflo r11
		//divu r1 / r9 (un)
		instmem [14] = 32'h0029001B;  //000000 00001 01001 00000 00000 011011  //divu r1 r9
		//sub r10 - r9 = -32(r12)
		instmem [15] = 32'h01496022;  //000000 01010 01001 01100 00000 100010  //sub r10 r9 r12
		//mult r6(40) * r12 (signed)
		instmem [16] = 32'h00CC0018;  //000000 00110 01100 00000 00000 011000  //mult r6 r12
		//div r6 / r12 (signed)
		instmem [17] = 32'h00CC001A;  //000000 00110 01100 00000 00000 011010  //div r6 r12
		//slt(12 11 13)
		instmem [18] = 32'h018B682A;  //000000 01100 01011 01101 00000 101010  //slt r12 r11 r13
		//slt(12 10 14)
		instmem [19] = 32'h018A702A;  //000000 01100 01010 01110 00000 101010  //slt r12 r10 r14
		//lui 15 -2
		instmem [20] = 32'h3C0FFFFF;  //001111 00000 01111 1111111111111111  //lui r15
 		//ori 15
		instmem [21] = 32'h35EFFFFE;  //001101 01111 01111 1111111111111110  //ori r15 r15 fffe
		//slt (12 15 16)
		instmem [22] = 32'h018F802A;  //000000 01100 01111 10000 00000 101010  //slt r12 r15 r16
		
		//mult r1 * r2
		instmem [23] = 32'h00220018;  //000000 00001 00010 00000 00000 011000  //mult r1 r2
    //mult r1 * r12
    instmem [24] = 32'h002C0018;  //000000 00001 01100 00000 00000 011000  //mult r1 r12
    //div r1 / r2
    instmem [25] = 32'h0022001A;  //000000 00001 00010 00000 00000 011010  //div r1 r2
    //div r12 / r6
    instmem [26] = 32'h0186001A;  //000000 01100 00110 00000 00000 011010  //div r12 r6
    //div r12 / r15
    instmem [27] = 32'h018F001A;  //000000 01100 01111 00000 00000 011010  //div r12 r15
    //sra 12 17
    instmem [28] = 32'h000C8883;  //000000 00000 01100 10001 00010 000011  //sra r12 r17

	 
      end
endmodule

